library verilog;
use verilog.vl_types.all;
entity mips32TOPTest2 is
end mips32TOPTest2;
