//------------------------------------------------------------------------------
//	Module:		Lab2Lock
//	Desc:			This module implements the functionality of a simple combination lock.
//					The lock uses 2 4-bit combination digits.
//					See the lab document for the suggested combination setting.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	Lab2Lock(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Enter,
			Digit,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			State,
			Open,
			Fail
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Parameters
	//--------------------------------------------------------------------------
	localparam	DIGIT_1	=	4'h2,
				DIGIT_2	=	4'h3,
				Locked = 3'b000, OK1 = 3'b001, Bad1 = 3'b010, Open1 = 3'b011, Bad2 = 3'b100;		
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Enter;
	input		[3:0]		Digit;
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output		[2:0]		State;
	output	reg				Open;
	output	reg				Fail;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	// place state encoding here
	
	//--------------------------------------------------------------------------
	 reg[2:0] state_on = Locked;
	assign State = state_on;
	 
	 	always @(state_on or Enter) begin
			case (state_on)

	 Locked: begin  //Locked

	 		Open = 1'b0;
			Fail = 1'b0;

	 end

	 OK1: begin //OK1
			Fail = 1'b0;
			Open = 1'b0;
	 end

	 Bad1: begin //BAD1
			Fail = 1'b1;
			Open = 1'b0;

	 end

	 Bad2: begin
			Fail = 1'b1;
			Open = 1'b0;
	 end

	Open1: begin
			Open = 1'b1;
			Fail = 1'b0;
	end	

	endcase

end
	
	always @ (posedge Clock, negedge Reset) begin
		
	

	if(~Reset)

	state_on <= Locked;
	else 
		case (state_on)

	 Locked: begin  //Locked
			
			if(Enter) begin
				if(Digit == DIGIT_1) state_on = OK1;
	 			else state_on <= Bad1;
			end

			else state_on <= Locked;
	 		
				 
				

	 end

	 OK1: begin //OK1

			if(Enter) begin
				if(Digit == DIGIT_2) state_on = Open1;
	 			else state_on <= Bad2;
			end

			else state_on <= OK1;

	 end

	 Bad1: begin //BAD1
			state_on <= Bad2;

	 end

	 Bad2: begin
			state_on <= Bad2;
	 end

	Open1: begin
			state_on <= Open1;
	end

	endcase

end


 
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------
	
	// Place you *fs Verilog here
	// You may find it useful to use a case statement to describe your FSM.

	//--------------------------------------------------------------------------
endmodule
//------------------------------------------------------------------------------
