library verilog;
use verilog.vl_types.all;
entity unitControlTb is
end unitControlTb;
