/***************************************************
 * Module: shiftLeft
 * Project: mips32
 * Description: Desloca 2 bits a esquerda (operação lógica)
 ***************************************************/
module shiftLeft(in, out);
	assign out = in << 2 ;
endmodule