// Universidade Estadual de Feira de Santana 
// TEC499 - MI - Sistemas Digitais
// Lab 3, 2016.1
//
// Module: ALU.v
// Desc:   32-bit ALU for the MIPS150 Processor
// Inputs: 
// 	A: 32-bit value
// 	B: 32-bit value
// 	ALUop: Selects the ALU's operation 
// 						
// Outputs:
// 	Out: The chosen function mapped to A and B.

`include "Opcode.vh"
`include "ALUop.vh"

module ALU(
    input [31:0] A,B,
    input [3:0] ALUop,
    output reg [31:0] Out
);
	
   wire signed [31:0] A_signed, B_signed;
	wire signed_comp;
	wire unsigned_comp;

  always@(*) begin 
  		

  		case(ALUop)

  			`ALU_ADDU: Out = A + B;
			`ALU_SUBU: Out = A - B;
			`ALU_SLT:  begin
							if(signed_comp == 1) Out = 32'd1;
							else Out = 32'd0;
				
						end
			`ALU_SLTU: begin
							if(unsigned_comp == 1) Out = 32'd1;
							else Out = 32'd0;
				
						end
			`ALU_AND: Out = A & B;
			`ALU_OR: Out = A | B;		
			`ALU_XOR: Out = A ^ B;
			`ALU_LUI: Out = B << 5'b10000;
			`ALU_SLLV: Out = B << A[4:0];
			`ALU_SRLV: Out = B >> A[4:0];
			`ALU_SRAV: Out = B_signed >>> A[4:0];
			`ALU_NOR: Out = (~A) & (~B);
			`ALU_XXX:  Out = 32'd0;



  		default: Out = 32'd0;

  		endcase
  end
  
  	
	assign signed_comp = ($signed(A) < $signed(B));
	assign unsigned_comp = A < B;
	assign B_signed = $signed(B);
  
endmodule
