`ifndef ALUOP
`define ALUOP

`define ALU_ADD  5'd0
`define ALU_DIV  5'd1
`define ALU_MUL  5'd2
`define ALU_SLT  5'd3
`define ALU_MFHI 5'd4
`define ALU_SUB  5'd5
`define ALU_XXX  5'd15

`endif //ALUOP
