/*************************************************************
 * Module: ulaControl
 * Project: mips32
 * Description: Só pra compilar o top
 ************************************************************/
module aluControl (opcode, funct, aluControlOut);
	input[5:0] opcode, funct;
	output[5:0] aluControlOut;

endmodule