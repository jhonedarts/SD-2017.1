library verilog;
use verilog.vl_types.all;
entity unitControlTest is
end unitControlTest;
